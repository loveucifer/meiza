# Op-Amp Non-Inverting Amplifier
# Basic non-inverting amplifier configuration

VIN dc_voltage 1V (0, -20) text="Input Signal"
U1 op_amp (50, 0) text="Operational Amplifier"
R1 resistor 1k (100, -30) text="Feedback Resistor"
R2 resistor 1k (100, 30) text="Ground Resistor"
VOUT test_point (150, 0) text="Amplified Output"
VCC dc_voltage 15V (0, -60) text="Positive Supply"
VEE dc_voltage -15V (0, 60) text="Negative Supply"
GND signal_ground (100, 80) text="Ground"

# Connections
VIN.+ -> U1.+  # Non-inverting input
U1.OUT -> R1.1  # Feedback to inverting input
R1.2 -> U1.-  # Connect to inverting input
R2.1 -> U1.-  # Connect to inverting input
R2.2 -> GND.GND
VCC.+ -> U1.V+  # Positive supply
VEE.- -> U1.V-  # Negative supply
VCC.- -> VEE.+  # Connect supplies together
VCC.- -> GND.GND
U1.OUT -> VOUT.TP  # Output