# RC Low-pass Filter
# This circuit implements a basic RC low-pass filter

VIN ac_voltage 1V (0, 0) text="Input Signal"
R1 resistor 1k (50, 0) text="Resistor"
C1 capacitor 10uF (100, 0) text="Filter Capacitor"
VOUT test_point (150, 0) text="Output"

GND signal_ground (75, 50) text="Circuit Ground"

# Connections
VIN.+ -> R1.1
R1.2 -> C1.1
C1.2 -> GND.GND
R1.2 -> VOUT.TP  # Output tap
VIN.- -> GND.GND