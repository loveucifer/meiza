# 555 Timer Astable Multivibrator
# This circuit creates an oscillator using a 555 timer

U1 timer_555 (0, 0) text="555 Timer"
R1 resistor 10k (50, -40) text="Timing Resistor 1"
R2 resistor 10k (50, 40) text="Timing Resistor 2"
C1 capacitor 10uF (100, 40) text="Timing Capacitor"
D1 diode (75, -40) text="Discharge Diode (optional)"
VCC dc_voltage 9V (0, -50) text="Supply"
GND signal_ground (100, 100) text="Ground"
OUT test_point (50, -80) text="Output"

# Connections
VCC.+ -> U1.VCC
U1.GND -> GND.GND
VCC.- -> GND.GND
U1.TRIG -> U1.THRES
U1.TRIG -> C1.1
C1.2 -> GND.GND
U1.DIS -> R2.1
R2.2 -> U1.THRES
R1.1 -> VCC.+
R1.2 -> U1.RESET
R1.2 -> U1.CONTROL
U1.OUT -> OUT.TP
D1.A -> R2.1
D1.K -> R1.2